0000000000011111111111 0000000000000000000000 0000000000011111111111 000
1111111111100000000000 0000000000000000000000 1111111111100000000000 010
0000000000000000000000 0000000000011111111111 0000000000011111111111 100
0000000000000000000000 1111111111100000000000 1111111111100000000000 110