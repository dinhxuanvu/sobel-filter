-------------------------------------------------------------------------------
-- File: memory_tb.vhd
-- Entity: memory_tb
-- Architecture: Behavioral
-- Author: Vu Dinh
-- Created: 12/03/2014
-- VHDL'93
-- Description: The following is the entity and architecture of a testbench
-- for memory module
-------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use IEEE.STD_LOGIC_TEXTIO.ALL;
use STD.TEXTIO.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all;

entity memory_tb is
end memory_tb;

architecture behavioral of memory_tb is

component memory is
  port
  (
    i_reset       :    in  std_logic;
    i_enable      :    in  std_logic;
    i_clock       :    in  std_logic;
    i_pixel       :    in  std_logic_vector(7 downto 0);
    o_ct          :    out std_logic_vector(71 downto 0)
  );
end component;

constant  period  :    time := 50 ns;
constant  delay   :    time := 10 ns;

signal s_i_reset  :    std_logic;
signal s_i_enable :    std_logic;
signal s_clk      :    std_logic;
signal s_i_pixel  :    std_logic_vector(7 downto 0);
signal s_o_ct     :    std_logic_vector(71 downto 0);

signal s_count    :    std_logic_vector(3 downto 0);
file INFILE: TEXT open READ_MODE is "memory_data";
-- pixel[7:0]     convolution table[71:0]
---  XXXXXXXX XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX 

begin
UUT: memory port map (s_i_reset, s_i_enable, s_clk, s_i_pixel, s_o_ct);
  
  verify : process
  
  variable    v_line       :   line; -- pointer to string
  variable    v_i_pixel    :   STD_LOGIC_VECTOR(7 DOWNTO 0);
  variable    v_o_ct       :   STD_LOGIC_VECTOR(71 DOWNTO 0);
  begin
    wait for DELAY;
    s_i_reset <= '1';
    wait until falling_edge(s_clk);
    s_i_reset <= '0';
    while not( endfile(INFILE)) loop  -- While not end of file,
      readline(INFILE, v_line);       -- read line of a file.
      read(v_line, v_i_pixel);    -- Each READ procedure extracts data
      read(v_line, v_o_ct);       -- from the beginning of the string
                                  -- value designed by parameter v_line.
      s_i_enable   <= '1';
      s_i_pixel    <= v_i_pixel;
      wait for DELAY;
      assert( v_o_ct=s_o_ct )
        report "convolution table is not correct";
      wait until rising_edge(s_clk);-- s_clk'EVENT;
    end loop;
    assert false
      report "done";
    wait;
  end process verify;

clock : process
begin
  s_clk <= '0';
  wait for period/2;
  s_clk <= '1';
  wait for period/2;
end process;
  		
end behavioral;