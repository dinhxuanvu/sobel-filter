-------------------------------------------------------------------------------
-- File: comparator.vhd
-- Entity: comparator
-- Architecture: Behavioral
-- Author: Drew Carlstedt, Vu Dinh
-- Created: 11/20/2014
-- VHDL'93
-- Description: The following is the entity and architecture of a 11-bit
-- comparator
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all;

entity comparator is
  port
  (
    i_enable     :    in  std_logic;
    i_d_n_e      :    in  std_logic_vector(21 downto 0);
    i_d_ne_nw    :    in  std_logic_vector(21 downto 0);
    o_d          :    out std_logic_vector(21 downto 0);
    o_dir        :    out std_logic_vector(2 downto 0)
  );
end comparator;

-------------------------------------------------------------------------------

architecture behavioral of comparator is

begin
  
  compare: process(i_d_n_e, i_d_ne_nw)
  variable v_d_n, v_d_e, v_d_ne, v_d_nw : std_logic_vector(10 downto 0);
  variable d_n_e, d_ne_nw               : std_logic_vector(10 downto 0);
  variable d_max                        : std_logic_vector(10 downto 0);
  variable dir_n_e, dir_ne_nw, dir_max  : std_logic_vector(2 downto 0);
  
  begin
    
    v_d_n   := i_d_n_e(21 downto 11);
    v_d_e   := i_d_n_e(10 downto 0);
    v_d_ne  := i_d_ne_nw(21 downto 11);
    v_d_nw  := i_d_ne_nw(10 downto 0);
    
    -- compare N and E
    if (abs(signed(v_d_n)) < abs(signed(v_d_e))) then
      d_n_e    := v_d_e;
      dir_n_e  := "000";
    else
      d_n_e    := v_d_n;
      dir_n_e  := "010";
    end if;
    -- compare NE and NW
    if (abs(signed(v_d_ne)) < abs(signed(v_d_nw))) then
      d_ne_nw   := v_d_nw;
      dir_ne_nw := "100";
    else
      d_ne_nw   := v_d_ne;
      dir_ne_nw := "110";
    end if;
    -- compare N/E and NE/NW
    if (abs(signed(d_n_e)) < abs(signed(d_ne_nw))) then
      d_max   := d_ne_nw;
      dir_max := dir_ne_nw;
    else
      d_max   := d_n_e;
      dir_max := dir_n_e;
    end if;
    
    -- if negative, opposite direction
    if (signed(d_max) < 0) then
      case dir_max is 
        when "010"  => -- N
              o_dir <= "011"; -- S
        when "000"  => -- E
              o_dir <= "001"; -- W
        when "110"  => -- NE
              o_dir <= "111"; -- SW
        when others => -- NW
              o_dir <= "101"; -- SE
      end case;
    else
      o_dir <= dir_max;
    end if;
    
    -- concatenate max derivative and perpendicular
    case dir_max is 
      when "010"  => -- N
            o_d   <= (d_max & v_d_e); 
      when "000"  => -- E
            o_d   <= (d_max & v_d_n);
      when "110"  => -- NE
            o_d   <= (d_max & v_d_nw);
      when others => -- NW
            o_d   <= (d_max & v_d_ne);
    end case;
  
  end process compare;
  
end behavioral;